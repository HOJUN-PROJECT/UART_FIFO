module clk_div_1khz_humid (
    input  clk,
    input  reset,
    output o_clk_1khz
);
    localparam DIV = 100000; // 100MHz / 100,000 = 1kHz

    reg [$clog2(DIV)-1:0] r_counter;
    reg r_clk_1khz;

    assign o_clk_1khz = r_clk_1khz;

    always @(posedge clk, posedge reset) begin
        if (reset) begin
            r_counter  <= 0;
            r_clk_1khz <= 1'b0;
        end else begin
            if (r_counter == DIV - 1) begin
                r_counter  <= 0;
                r_clk_1khz <= 1'b1;
            end else begin
                r_counter  <= r_counter + 1;
                r_clk_1khz <= 1'b0;
            end
        end
    end
endmodule
